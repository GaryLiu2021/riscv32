// tb
//`define ALL




`define     CLK_FRE             50 // MHz

// AHB
`define     AHB_ADDR_WIDTH      32
`define     AHB_DATA_WIDTH      32

// UART
`define     BAUD_RATE           115200

// ram
`define     RAM_DEPTH           65536
    //实际上该是65536